/*
 * First module.
 *  dependencies:
 *	initial procedural block
 *	sequential block
 */

module main;

	initial
		begin
		end

endmodule
